 .option post
Vin	1	0	SIN	0V 1V 10meg
R1	1	2	2k
C1	2	0	1p
L1	2	3	1n
R2	3	0	3k
.tran 1ns 1us
.end