.option post
V1	1	0	5V
R1	1	2	330
D1	2	0	diode
.model	diode	D
.tran	0.1ns	1ns
.end