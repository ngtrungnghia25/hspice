.option post
V1	0	1	5V
D1	0	1	mod1
.model	mod1	d
.tran	0.1ns	1ns
.end